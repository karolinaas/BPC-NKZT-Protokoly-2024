** Profile: "SCHEMATIC1-AC char"  [ D:\student\247759\Zesilovac AC char\zesilovac ac char-schematic1-ac char.sim ] 

** Creating circuit file "zesilovac ac char-schematic1-ac char.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "C:\Program Files\Orcad\PSpice\UserLib\Tube_IM.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\zesilovac ac char-SCHEMATIC1.net" 


.END
