** Profile: "SCHEMATIC1-Prevodni char"  [ D:\student\247759\Prevodni char\prevodni char-schematic1-prevodni char.sim ] 

** Creating circuit file "prevodni char-schematic1-prevodni char.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "C:\Program Files\Orcad\PSpice\UserLib\Tube_IM.lib" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 -3 0 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\prevodni char-SCHEMATIC1.net" 


.END
